`ifndef ULTRA_CORE_ENV_PKG__SV
`define ULTRA_CORE_ENV_PKG__SV

  package ultra_core_env_pkg;

    // Import UVM
    import uvm_pkg::*;
    import ultra_core_seq_pkg::*;
    import ultra_core_regs_pkg::*;
    import ultra_core_agent_pkg::*;
    `include "uvm_macros.svh"

    // Import UVM
    `include "ultra_core_sb.sv"
    `include "ultra_core_cov.sv"
    `include "ultra_core_env.sv"
  endpackage

`endif

//End of ultra_core_env_pkg
