`ifndef ULTRA_CORE_REGS_PKG__SV
`define ULTRA_CORE_REGS_PKG__SV

  package ultra_core_regs_pkg;

    // Import UVM
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Include Reg Model UVCs

  endpackage

`endif

//End of ultra_core_regs_pkg
